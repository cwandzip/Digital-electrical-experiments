module data2ascii (code, ascii);
	input [7:0] code;
	output [7:0] ascii;
/* verilator lint_off WIDTHEXPAND */
	MuxKeyWithDefault #(36, 8, 8) mux0 (ascii, code, 8'b00000000, {
		//数字
		8'h16, 8'b00110001, //1
		8'h1E, 8'b00110010, 
		8'h26, 8'b00110011, 
		8'h25, 8'b00110100, 
		8'h2E, 8'b00110101, 
		8'h36, 8'b00110110, 
		8'h3D, 8'b00110111, 
		8'h3E, 8'b00111000, 
		8'h46, 8'b00111001, 
		8'h45, 8'b00110000, //0
		//字母
		8'h1C, 8'b01100001, //a
		8'h32, 8'b01100010, //b
		8'h21, 8'b01100011, 
		8'h23, 8'b01100100, 
		8'h24, 8'b01100101, 
		8'h2B, 8'b01100110, 
		8'h34, 8'b01100111, 
		8'h33, 8'b01101000, 
		8'h43, 8'b01101001, 
		8'h3B, 8'b01101010, 
		8'h42, 8'b01101011, 
		8'h4B, 8'b01101100, 
		8'h3A, 8'b01101101, 
		8'h31, 8'b01101110, 
		8'h44, 8'b01101111, 
		8'h4D, 8'b01110000, 
		8'h15, 8'b01110001, 
		8'h2D, 8'b01110010, 
		8'h1B, 8'b01110011, 
		8'h2C, 8'b01110100, 
		8'h3C, 8'b01110101, 
		8'h2A, 8'b01110110, 
		8'h1D, 8'b01110111, 
		8'h22, 8'b01111000, 
		8'h35, 8'b01111001, 
		8'h1A, 8'b01111010
	});
/* verilator lint_off WIDTHEXPAND */
endmodule
